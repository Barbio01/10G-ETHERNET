-- EMACS settings: -*- tab-width: 2; indent-tabs-mode: nil -*-
-- vim: tabstop=2:shiftwidth=2:expandtab
-- kate: tab-width 2; replace-tabs on; indent-width 2;

------------------------------<-    80 chars    ->------------------------------
--! @file
--! @brief Interfaces context of the project
--! @details Contains the full list of interfaces,
--! inherits from constants.vhd.
--! @author Steffen Stärz <steffen.staerz@cern.ch>
--------------------------------------------------------------------------------

--! @cond
context interfaces is

  library IEEE;
      use IEEE.STD_LOGIC_1164.ALL;  -- Defines std_logic and std_logic_vector
      use IEEE.NUMERIC_STD.ALL;

  library PoC;
    use PoC.utils.all;

  library fpga;
    --context fpga.constants;
    use fpga.fpga_if.all;

end context interfaces;

--! @endcond
